module torri

pub fn encode_jpeg(file_path string) []byte {
	return 'Ok'.bytes()
}

